localparam W_BYTES = 103636;
localparam X_BYTES = 648;
localparam Y_BYTES = 73736;
localparam X_BYTES_ALL = 105008;
