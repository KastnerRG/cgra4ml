localparam N_BUNDLES = 6;

Bundle_t bundles [N_BUNDLES] = '{
  '{ w_wpt:2368,  w_wpt_p0:2368,  x_wpt:424,  x_wpt_p0:424,  y_wpt:16,  y_wpt_last:96,  y_nl:4,  y_w:3,  n_it:8,  n_p:3 },
  '{ w_wpt:2208,  w_wpt_p0:2208,  x_wpt:840,  x_wpt_p0:840,  y_wpt:24,  y_wpt_last:96,  y_nl:4,  y_w:5,  n_it:6,  n_p:8 },
  '{ w_wpt:1568,  w_wpt_p0:608,  x_wpt:1256,  x_wpt_p0:424,  y_wpt:32,  y_wpt_last:96,  y_nl:4,  y_w:6,  n_it:4,  n_p:6 },
  '{ w_wpt:1176,  w_wpt_p0:312,  x_wpt:2088,  x_wpt_p0:424,  y_wpt:64,  y_wpt_last:128,  y_nl:4,  y_w:7,  n_it:3,  n_p:4 },
  '{ w_wpt:1176,  w_wpt_p0:744,  x_wpt:6248,  x_wpt_p0:3752,  y_wpt:192,  y_wpt_last:192,  y_nl:4,  y_w:8,  n_it:3,  n_p:2 },
  '{ w_wpt:392,  w_wpt_p0:272,  x_wpt:398,  x_wpt_p0:268,  y_wpt:192,  y_wpt_last:192,  y_nl:2,  y_w:1,  n_it:1,  n_p:427 }
};