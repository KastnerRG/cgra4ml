`define VALID_PROB 1000 
`define READY_PROB 1000