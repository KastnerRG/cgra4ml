localparam W_BYTES = 206240;
localparam X_BYTES = 1272;
localparam X_BYTES_ALL = 201200;
