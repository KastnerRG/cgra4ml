
`define VALID_PROB 1000 
`define READY_PROB 1000 
`define CLK_PERIOD 4.0 
`define INPUT_DELAY_NS  0.8ns
`define OUTPUT_DELAY_NS 0.8ns
