
`define VALID_PROB 1000 
`define READY_PROB 1000 
`define CLK_PERIOD 6.7 
`define INPUT_DELAY_NS  1.3ns
`define OUTPUT_DELAY_NS 1.3ns
