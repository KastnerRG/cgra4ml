`define VALID_PROB 1 
`define READY_PROB 100