`define VALID_PROB 100 
`define READY_PROB 100