
`define VALID_PROB 10 
`define READY_PROB 100 
`define CLK_PERIOD 6.7 
`define INPUT_DELAY_NS  1.3ns
`define OUTPUT_DELAY_NS 1.3ns
