`define VALID_PROB 10 
`define READY_PROB 100