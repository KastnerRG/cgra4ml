
`define VALID_PROB 100 
`define READY_PROB 10 
`define CLK_PERIOD 4.0 
`define INPUT_DELAY_NS  0.8ns
`define OUTPUT_DELAY_NS 0.8ns
